`include "eth_axis_rx_module.sv";
`include "eth_axis_tx_module.sv";
`include "eth_mac_10g.sv";
`include "eth_phy_10g.sv";
module eth_axi_stream_top #
(

parameter DATA_WIDTH = 64,

parameter HDR_WIDTH = 2,

parameter KEEP_WIDTH = (DATA_WIDTH/8),

parameter CTRL_WIDTH = (DATA_WIDTH/8),

parameter ENABLE_PADDING = 1,

parameter ENABLE_DIC = 1,

parameter MIN_FRAME_LENGTH = 64,

parameter PTP_TS_ENABLE = 0,

parameter PTP_TS_FMT_TOD = 1,

parameter PTP_TS_WIDTH = PTP_TS_FMT_TOD ? 96 : 64,

parameter TX_PTP_TS_CTRL_IN_TUSER = 0,

parameter TX_PTP_TAG_ENABLE = PTP_TS_ENABLE,

parameter TX_PTP_TAG_WIDTH = 16,

parameter TX_USER_WIDTH = (PTP_TS_ENABLE ? (TX_PTP_TAG_ENABLE ? TX_PTP_TAG_WIDTH : 0) + (TX_PTP_TS_CTRL_IN_TUSER ? 1 : 0) : 0) + 1,

parameter RX_USER_WIDTH = (PTP_TS_ENABLE ? PTP_TS_WIDTH : 0) + 1,

parameter PFC_ENABLE = 0,

parameter PAUSE_ENABLE = PFC_ENABLE

)
(
  input wire rx_clk,
  input wire rx_rst,
  input wire tx_clk,
  input wire tx_rst,
  input wire [DATA_WIDTH-1:0]tx_axis_tdata,
  input wire [KEEP_WIDTH-1:0]tx_axis_tkeep,
  input wire tx_axis_tvalid, 
  input wire tx_axis_tready, 
  input wire tx_axis_tlast,
  input wire [TX_USER_WIDTH-1:0] tx_axis_tuser,
  output wire [DATA_WIDTH-1:0] rx_axis_tdata,
  output wire [KEEP_WIDTH-1:0] rx_axis_tkeep,
  output wire rx_axis_tvalid,
  output wire rx_axis_tlast,
  output wire [RX_USER_WIDTH-1:0] rx_axis_tuser,
  input  wire  [DATA_WIDTH-1:0]  xgmii_rxd,
  input  wire  [CTRL_WIDTH-1:0]  xgmii_rxc,
  output wire  [DATA_WIDTH-1:0]  xgmii_txd,
  output wire  [CTRL_WIDTH-1:0]  xgmii_txc,
  input  wire [PTP_TS_WIDTH-1:0] tx_ptp_ts,
  input  wire [PTP_TS_WIDTH-1:0] rx_ptp_ts,
  output wire [PTP_TS_WIDTH-1:0] tx_axis_ptp_ts,
  output wire [PTP_TS_WIDTH-1:0] tx_axis_ptp_ts_tag,
  output wire tx_axis_ptp_ts_valid, 
  input wire tx_lfc_req,
  input wire tx_lfc_resend,
  input wire rx_lfc_en,
  input wire rx_lfc_req,
  input wire rx_lfc_ack, 
  input wire [7:0] tx_pfc_req,
  input wire tx_pfc_resend,
  input wire [7:0] rx_pfc_en,
  input wire [7:0] rx_pfc_req,
  input wire [7:0] rx_pfc_ack,
//*Pause Interface
  input wire tx_lfc_pasue_en,
  input wire tx_pause_req,
  output wire tx_pause_ack,
/* status */ 
 output wire [1:0] tx_start_packet,
 output wire tx_error_underflow,
 output wire [1:0] rx_start_packet,
 output wire rx_error_bad_frame,
 output wire rx_error_bad_fcs,
 output wire stat_tx_mcf,
 output wire stat_rx_mcf,
 output wire stat_tx_lfc_pkt,
 output wire stat_tx_lfc_xon,
 output wire stat_tx_lfc_xoff,
 output wire stat_tx_lfc_paused,
 output wire stat_tx_pfc_pkt,
 output wire stat_tx_pfc_xon,
 output wire stat_tx_pfc_xoff,
 output wire stat_tx_pfc_paused,
 output wire stat_rx_lfc_pkt,
 output wire stat_rx_lfc_xon,
 output wire stat_rx_lfc_xoff,
 output wire stat_rx_lfc_paused,
 output wire stat_rx_pfc_pkt,
 output wire stat_rx_pfc_xon,
 output wire stat_rx_pfc_xoff,
 output wire stat_rx_pfc_paused,
/*
*Configuration
*/
input wire [7:0] cfg_ifg,
input wire cfg_tx_enable,
input wire cfg_rx_enable,
input wire [47:0]  cfg_mcf_rx_eth_dst_mcast,
input wire  cfg_mcf_rx_check_eth_dst_mcast,
input wire [47:0] cfg_mcf_rx_eth_dst_ucast,
input wire cfg_mcf_rx_check_eth_dst_ucast,
input wire [47:0] cfg_mcf_rx_eth_src,
input wire cfg_mcf_rx_check_eth_src,
input wire [15:0] cfg_mcf_rx_eth_type,
input wire [15:0] cfg_mcf_rx_opcode_lfc,
input wire cfg_mcf_rx_check_opcode_lfc,
input wire [15:0] cfg_mcf_rx_opcode_pfc,
input wire cfg_mcf_rx_check_opcode_pfc,
input wire cfg_mcf_rx_forward,
input wire cfg_mcf_rx_enable,
input wire [47:0] cfg_tx_lfc_eth_dst,
input wire [47:0] cfg_tx_lfc_eth_src,
input wire [15:0] cfg_tx_lfc_eth_type,
input wire [15:0] cfg_tx_lfc_opcode,
input wire cfg_tx_lfc_en,
input wire [15:0] cfg_tx_lfc_quanta,
input wire [15:0] cfg_tx_lfc_refresh,
input wire [47:0] cfg_tx_pfc_eth_dst,
input wire [47:0] cfg_tx_pfc_eth_src,
input wire [15:0] cfg_tx_pfc_eth_type,
input wire [15:0] cfg_tx_pfc_opcode,
input wire cfg_tx_pfc_en,
input wire [8*16-1:0] cfg_tx_pfc_quanta,
input wire [8*16-1:0] cfg_tx_pfc_refresh,
input wire [15:0] cfg_rx_lfc_opcode,
input wire cfg_rx_lfc_en,
input wire [15:0] cfg_rx_pfc_opcode,
input wire cfg_rx_pfc_en, 

/*
* XGMII interface
*/

//input wire [DATA_WIDTH-1:0] xgmii_txd,
//input wire [CTRL_WIDTH-1:0] xgmii_txc,
//output wire [DATA_WIDTH-1:0] xgmii_rxd,
//output wire [CTRL_WIDTH-1:0] xgmii_rxc,

/*
* SERDES interface
*/

output wire [DATA_WIDTH-1:0] serdes_tx_data,
output wire [HDR_WIDTH-1:0] serdes_tx_hdr,
input wire [DATA_WIDTH-1:0] serdes_rx_data,
input wire [HDR_WIDTH-1:0] serdes_rx_hdr,
output wire serdes_rx_bitslip,
output wire serdes_rx_reset_req,

/*
* Status
*/

output wire tx_bad_block,
output wire [6:0] rx_error_count,
output wire rx_bad_block,
output wire rx_sequence_error,
output wire rx_block_lock,
output wire rx_high_ber,
output wire rx_status,

/*
* Configuration
*/

input wire cfg_tx_prbs31_enable,
input wire cfg_rx_prbs31_enable

);

wire [DATA_WIDTH-1:0] top_rx_axis_tdata;
wire [KEEP_WIDTH-1:0] top_rx_axis_tkeep;
wire top_rx_axis_tvalid;
wire top_rx_axis_tlast;
wire [RX_USER_WIDTH-1:0] top_rx_axis_tuser;

wire [DATA_WIDTH-1:0]top_tx_axis_tdata;
wire [KEEP_WIDTH-1:0]top_tx_axis_tkeep;
wire top_tx_axis_tvalid;
wire top_tx_axis_tready;
wire top_tx_axis_tlast;
wire [TX_USER_WIDTH-1:0] tx_axis_tuser;


wire [7:0] top_cfg_ifg;
wire cfg_tx_enable;
wire cfg_rx_enable;
wire cfg_mcf_rx_eth_dst_mcast;
wire cfg_mcf_rx_check_eth_dst_mcast;
wire cfg_mcf_rx_eth_dst_ucast;
wire cfg_mcf_rx_check_eth_dst_ucast;
wire cfg_mcf_rx_eth_src;
wire cfg_mcf_rx_check_eth_src;
wire cfg_mcf_rx_eth_type;
wire cfg_mcf_rx_opcode_lfc;
wire cfg_mcf_rx_opcode_pfc;
wire cfg_mcf_rx_check_opcode_pfc;
wire cfg_mcf_rx_forward;
wire cfg_mcf_rx_enable;
wire cfg_tx_lfc_eth_dst;
wire cfg_tx_lfc_eth_src;
wire cfg_tx_lfc_eth_type;
wire cfg_tx_lfc_opcode;
wire cfg_tx_lfc_en;
wire cfg_tx_lfc_quanta;
wire cfg_tx_lfc_refresh;
wire cfg_tx_pfc_eth_dst;
wire cfg_tx_pfc_eth_src;
wire cfg_tx_pfc_eth_type;
wire cfg_tx_pfc_opcode;
wire cfg_tx_pfc_en;
wire cfg_tx_pfc_quanta;
wire cfg_tx_pfc_refresh;
wire cfg_rx_lfc_opcode;
wire cfg_rx_lfc_en;
wire cfg_rx_pfc_opcode;
wire cfg_rx_pfc_en;

wire [PTP_TS_WIDTH-1:0] top_tx_ptp_ts;
wire [PTP_TS_WIDTH-1:0] top_rx_ptp_ts;
wire [PTP_TS_WIDTH-1:0] top_tx_axis_ptp_ts;
wire [PTP_TS_WIDTH-1:0] top_tx_axis_ptp_ts_tag;
wire  top_tx_axis_ptp_ts_valid;

//Link Flow control
wire top_tx_lfc_req;
wire top_tx_lfc_resend;
wire top_rx_lfc_en;
wire top_rx_lfc_req;
wire top_rx_lfc_ack;

   
wire [7:0] top_tx_pfc_req;
wire top_tx_pfc_resend;
wire [7:0] top_rx_pfc_en;
wire [7:0] top_rx_pfc_req;
wire [7:0] top_rx_pfc_ack;

wire top_tx_lfc_pause_en;
wire top_tx_pause_req;
wire top_tx_pause_ack;

//phy signals
wire rx_clk;
wire rx_rst;
wire tx_clk;
wire tx_rst;

wire top_xgmii_txd;
wire top_xgmii_txc;
wire top_xgmii_rxd;
wire top_xgmii_rxc;

wire serdes_tx_data;
wire serdes_tx_hdr;
wire serdes_rx_data;
wire serdes_rx_hdr;
wire serdes_rx_bitslip;
wire serdes_rx_reset_req;

wire tx_bad_block;
wire [6:0] rx_error_count;
wire rx_bad_clock;
wire rx_sequence_error;
wire rx_block_lock;
wire rx_high_ber;
wire rx_status;

wire cfg_tx_prbs31_enable;
wire cfg_rx_prbs31_enable;

wire top_rx_clk;
wire top_rx_rst;
wire top_tx_clk;
wire top_tx_rst;

wire [1:0] top_tx_start_packet;
wire top_tx_error_underflow;
wire [1:0] top_rx_start_packet;
wire top_rx_error_bad_frame;
wire top_rx_error_bad_fcs;
wire top_sta_tx_mcf;
wire top_stat_tx_mcf;
wire top_stat_tx_lfc_pkt;
wire top_stat_tx_lfc_xon;
wire top_stat_tx_lfc_xoff;
wire top_stat_tx_lfc_paused;
wire top_stat_tx_pfc_pkt;
wire [7:0] top_stat_tx_pfc_xon;
wire [7:0] top_stat_tx_pfc_xoff;
wire [7:0] top_stat_tx_pfc_paused;

wire top_stat_rx_lfc_pkt;
wire top_stat_rx_lfc_xon;
wire top_stat_rx_lfc_xoff;
wire top_stat_rx_lfc_paused;
wire top_stat_rx_pfc_pkt;
wire [7:0] top_stat_rx_pfc_xon;
wire [7:0] top_stat_rx_pfc_xoff;
wire [7:0] top_stat_rx_pfc_paused;

wire [7:0] top_cfg_ifg;
wire top_cfg_tx_enable;
wire top_cfg_rx_enable;
wire [47:0]  top_cfg_mcf_rx_eth_dst_mcast;
wire  top_cfg_mcf_rx_check_eth_dst_mcast;
wire [47:0] top_cfg_mcf_rx_eth_dst_ucast;
wire top_cfg_mcf_rx_check_eth_dst_ucast;
wire [47:0] top_cfg_mcf_rx_eth_src;
wire top_cfg_mcf_rx_check_eth_src;
wire [15:0] top_cfg_mcf_rx_eth_type;
wire [15:0] top_cfg_mcf_rx_opcode_lfc;
wire top_cfg_mcf_rx_check_opcode_lfc;
wire [15:0] top_cfg_mcf_rx_opcode_pfc;
wire top_cfg_mcf_rx_check_opcode_pfc;
wire top_cfg_mcf_rx_forward;
wire top_cfg_mcf_rx_enable;
wire [47:0] top_cfg_tx_lfc_eth_dst;
wire [47:0] top_cfg_tx_lfc_eth_src;
wire [15:0] top_cfg_tx_lfc_eth_type;
wire [15:0] top_cfg_tx_lfc_opcode;
wire top_cfg_tx_lfc_en;
wire [15:0] top_cfg_tx_lfc_quanta;
wire [15:0] top_cfg_tx_lfc_refresh;
wire [47:0] top_cfg_tx_pfc_eth_dst;
wire [47:0] top_cfg_tx_pfc_eth_src;
wire [15:0] top_cfg_tx_pfc_eth_type;
wire [15:0] top_cfg_tx_pfc_opcode;
wire top_cfg_tx_pfc_en;
wire [8*16-1:0] top_cfg_tx_pfc_quanta;
wire [8*16-1:0] top_cfg_tx_pfc_refresh;
wire [15:0] top_cfg_rx_lfc_opcode;
wire top_cfg_rx_lfc_en;
wire [15:0] top_cfg_rx_pfc_opcode;
wire top_cfg_rx_pfc_en;

eth_mac_10g  #(.DATA_WIDTH(DATA_WIDTH),

               .KEEP_WIDTH(DATA_WIDTH/8),

               .CTRL_WIDTH(DATA_WIDTH/8),

               .ENABLE_PADDING(1),

               .ENABLE_DIC(1),

               .MIN_FRAME_LENGTH(64),

               .PTP_TS_ENABLE(0),

               .PTP_TS_FMT_TOD(1),

               .PTP_TS_WIDTH(96),

               .TX_PTP_TS_CTRL_IN_TUSER(0),

               .TX_PTP_TAG_ENABLE(0),

               .TX_PTP_TAG_WIDTH(16),

               .TX_USER_WIDTH(1),

               .RX_USER_WIDTH(1),

               .PFC_ENABLE(0),

               .PAUSE_ENABLE(0)

)

eth_mac_10g_inst ( 
 .rx_clk(top_rx_clk),
 .rx_rst(top_rx_rst),
 .tx_clk(top_tx_clk),
 .tx_rst(top_tx_rst), 
  
  //AXI i/p
 .tx_axis_tdata(top_tx_axis_tdata),
 .tx_axis_tkeep(top_tx_axis_tkeep),
 .tx_axis_tvalid(top_axis_tvalid),
 .tx_axis_tready(top_axis_tready),
 .tx_axis_tlast(top_axis_tlast),
 .tx_axis_tuser(top_axis_tuser),

 //AXI o/p
  .rx_axis_tdata(top_rx_axis_tdata),
  .rx_axis_tkeep(top_rx_axis_tkeep),
  .rx_axis_tvalid(top_rx_axis_tvalid),
  .rx_axis_tlast(top_rx_axis_tlast),
  .rx_axis_tuser(top_rx_axis_tuser),

 //XGMII interface

  .xgmii_rxd(top_xgmii_rxd),
  .xgmii_rxc(top_xgmii_rxc),
  .xgmii_txd(top_xgmii_txd),
  .xgmii_txc(top_xgmii_txc),

  .tx_ptp_ts(top_tx_ptp_ts),
  .rx_ptp_ts(top_rx_ptp_ts),
  .tx_axis_ptp_ts(top_tx_axis_ptp_ts),
  .tx_axis_ptp_ts_tag(top_tx_axis_ptp_ts_tag),
  .tx_axis_ptp_ts_valid(top_tx_axis_ptp_ts_valid),

  .tx_lfc_req(top_tx_lfc_req),
  .tx_lfc_resend(top_tx_lfc_resend),
  .rx_lfc_en(top_rx_lfc_en),
  .rx_lfc_req(top_rx_lfc_req),
  .rx_lfc_ack(top_rx_lfc_ack), 

  .tx_pfc_req(top_tx_pfc_req),
  .tx_pfc_resend(top_tx_pfc_resend),
  .rx_pfc_en(top_rx_pfc_en),
  .rx_pfc_req(top_rx_pfc_req),
  .rx_pfc_ack(top_rx_pfc_ack),

  
  .tx_lfc_pause_en(top_tx_lfc_pause_en),
  .tx_pause_req(top_tx_pause_req),
  .tx_pause_ack(top_tx_pause_ack),
  
  .tx_start_packet(top_tx_start_packet),
  .tx_error_underflow(top_tx_error_underflow),
  .rx_start_packet(top_rx_start_packet),
  .rx_error_bad_frame(top_rx_error_bad_frame),
  .rx_error_bad_fcs(top_ex_error_bad_fcs),
  .stat_tx_mcf(top_stat_tx_mcf),
  .stat_rx_mcf(top_stat_rx_mcf),
  .stat_tx_lfc_pkt(top_stat_tx_lfc_pkt),
  .stat_tx_lfc_xon(top_stat_tx_lfc_xon),
  .stat_tx_lfc_xoff(top_stat_tx_lfc_xoff),
  .stat_tx_lfc_paused(top_stat_tx_lfc_paused),
  .stat_tx_pfc_pkt(top_stat_tx_pfc_pkt),
  .stat_tx_pfc_xon(top_stat_tx_pfc_xon),
  .stat_tx_pfc_xoff(top_stat_tx_pfc_xoff),
  .stat_tx_pfc_paused(top_stat_tx_pfc_pasued),
  .stat_rx_lfc_pkt(top_stat_rx_lfc_pkt),
  .stat_rx_lfc_xon(top_stat_rx_lfc_xon),
  .stat_rx_lfc_xoff(top_stat_rx_lfc_xoff),
  .stat_rx_lfc_paused(top_stat_rx_lfc_pasued),
  .stat_rx_pfc_pkt(top_stat_rx_pfc_pkt),
  .stat_rx_pfc_xon(top_stat_rx_pfc_xon),
  .stat_rx_pfc_xoff(top_stat_rx_pfc_xoff),
  .stat_rx_pfc_paused(top_stat_rx_pfc_paused),
/*
*Configuration
*/
 .cfg_ifg(top_cfg_ifg),
 .cfg_tx_enable(top_cfg_tx_enable),
 .cfg_rx_enable(top_cfg_rx_enable),
 .cfg_mcf_rx_eth_dst_mcast(top_cfg_mcf_rx_eth_dst_mcast),
 .cfg_mcf_rx_check_eth_dst_mcast(top_cfg_mcf_rx_check_eth_dst_mcast),
 .cfg_mcf_rx_eth_dst_ucast(top_cfg_mcf_rx_eth_dst_ucast),
 .cfg_mcf_rx_check_eth_dst_ucast(top_cfg_mcf_rx_check_eth_dst_ucast),
 .cfg_mcf_rx_eth_src(top_cfg_mcf_rx_eth_src),
 .cfg_mcf_rx_check_eth_src(top_cfg_mcf_rx_check_eth_src),
 .cfg_mcf_rx_eth_type(top_cfg_mcf_rx_eth_type),
 .cfg_mcf_rx_opcode_lfc(top_cfg_mcf_rx_opcode_lfc),
 .cfg_mcf_rx_check_opcode_lfc(top_cfg_mcf_rx_check_opcode_lfc),
 .cfg_mcf_rx_opcode_pfc(top_cfg_mcf_rx_opcode_pfc),
 .cfg_mcf_rx_check_opcode_pfc(top_cfg_mcf_rx_check_opcode_pfc),
 .cfg_mcf_rx_forward(top_cfg_mcf_rx_forward),
 .cfg_mcf_rx_enable(top_cfg_mcf_rx_enable),
 .cfg_tx_lfc_eth_dst(top_cfg_tx_lfc_eth_dst),
 .cfg_tx_lfc_eth_src(top_cfg_tx_lfc_eth_src),
 .cfg_tx_lfc_eth_type(top_cfg_tx_lfc_eth_type),
 .cfg_tx_lfc_opcode(top_cfg_tx_lfc_opcode),
 .cfg_tx_lfc_en(top_cfg_tx_lfc_en),
 .cfg_tx_lfc_quanta(top_cfg_tx_lfc_en),
 .cfg_tx_lfc_refresh(top_cfg_tx_lfc_refresh),
 .cfg_tx_pfc_eth_dst(top_cfg_tx_pfc_eth_dst),
 .cfg_tx_pfc_eth_src(top_cfg_tx_pfc_eth_dst),
 .cfg_tx_pfc_eth_type(top_cfg_tx_pfc_eth_type),
 .cfg_tx_pfc_opcode(top_cfg_tx_pfc_opcode),
 .cfg_tx_pfc_en(top_cfg_tx_pfc_en),
 .cfg_tx_pfc_quanta(top_cfg_tx_pfc_quanta),
 .cfg_tx_pfc_refresh(top_cfg_tx_pfc_refresh),
 .cfg_rx_lfc_opcode(top_cfg_rx_lfc_opcode),
 .cfg_rx_lfc_en(top_cfg_rx_lfc_en),
 .cfg_rx_pfc_opcode(top_cfg_rx_pfc_opcode),
 .cfg_rx_pfc_en(top_cfg_rx_pfc_en) 
); 

eth_phy_10g  #(

.DATA_WIDTH(DATA_WIDTH),
.CTRL_WIDTH(DATA_WIDTH/8),
.HDR_WIDTH(2),
.BIT_REVERSE(0),
.SCRAMBLER_DISABLE(0),
.PRBS31_ENABLE(0),
.TX_SERDES_PIPELINE(0),
.RX_SERDES_PIPELINE(0),
.BITSLIP_HIGH_CYCLES(1),
.BITSLIP_LOW_CYCLES(8),
.COUNT_125US(125000/6.4)
)
eth_phy_10g_inst ( 
   .rx_clk(top_rx_clk),
   .rx_rst(top_rx_rst),
   .tx_clk(top_tx_clk),
   .tx_rst(top_tx_rst),
   
   .xgmii_txd(top_xgmii_txd),
   .xgmii_txc(top_xgmii_txc),
   .xgmii_rxd(top_xgmii_rxd),
   .xgmii_rxc(top_xgmii_rxc),

   .serdes_tx_data(top_serdes_tx_data),
   .serdes_tx_hdr(top_serdes_tx_hdr),    
   .serdes_rx_data(top_serdes_rx_data),
   .serdes_rx_hdr(top_serdes_rx_hdr),
   .serdes_rx_bitslip(top_serdes_rx_bitslip),
   .serdes_rx_reset_req(top_serdes_rx_reset_req),
  
   .tx_bad_block(top_tx_bad_block),
   .rx_error_count(top_rx_error_count),
   .rx_bad_block(top_rx_bad_block),
   .rx_sequence_error(top_rx_sequence_error),
   .rx_block_lock(top_rx_block_lock),
   .rx_high_ber(top_rx_high_ber),
   .rx_status(top_rx_status),
   .cfg_tx_prbs31_enable(top_cfg_tx_prbs31_enable),
   .cfg_rx_prbs31_enable(top_cfg_rx_prbs31_enable)
   );
   
endmodule:eth_axi_stream_top
